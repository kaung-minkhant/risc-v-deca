LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY data_path IS
    PORT (
        -- reset and clock
        clk
    );
END data_path;

ARCHITECTURE rtl OF data_path IS

BEGIN

END ARCHITECTURE;